module Clock(CLOCK);
    output reg CLOCK;
initial begin
  #1	CLOCK = 1;
  #1	CLOCK = 0;
  #1	CLOCK = 1;
  #1	CLOCK = 0;
  #1	CLOCK = 1;
  #1	CLOCK = 0;
  #1	CLOCK = 1;
  #1	CLOCK = 0;
  #1	CLOCK = 1;
  #1	CLOCK = 0;
  #1	CLOCK = 1;
  #1	CLOCK = 0;
  #1	CLOCK = 1;
  #1	CLOCK = 0;
  #1	CLOCK = 1;
  #1	CLOCK = 0;
  #1	CLOCK = 1;
  #1	CLOCK = 0;
  #1	CLOCK = 1;
  #1	CLOCK = 0;
  #1	CLOCK = 1;
  #1	CLOCK = 0;
  #1	CLOCK = 1;
  #1	CLOCK = 0;
  #1	CLOCK = 1;
  #1	CLOCK = 0;
  #1	CLOCK = 1;
  #1	CLOCK = 0;
  #1	CLOCK = 1;
  #1	CLOCK = 0;
  #1	CLOCK = 1;
  #1	CLOCK = 0;
  #1	CLOCK = 1;
  #1	CLOCK = 0;
  #1	CLOCK = 1;
  #1	CLOCK = 0;
  #1	CLOCK = 1;
  #1	CLOCK = 0;
  #1	CLOCK = 1;
  #1	CLOCK = 0;
  #1	CLOCK = 1;
  #1	CLOCK = 0;
  #1	CLOCK = 1;
  #1	CLOCK = 0;
  #1	CLOCK = 1;
  #1	CLOCK = 0;
  #1	CLOCK = 1;
  #1	CLOCK = 0;
  #1	CLOCK = 1;
  #1	CLOCK = 0;
  #1	CLOCK = 1;
  #1	CLOCK = 0;
  #1	CLOCK = 1;
  #1	CLOCK = 0;
  #1	CLOCK = 1;
  #1	CLOCK = 0;
  #1	CLOCK = 1;
  #1	CLOCK = 0;
  #1	CLOCK = 1;
  #1	CLOCK = 0;

end


endmodule
